* ============================================================================
* RL Lowpass Filter — First-order
* PedalKernel Validation Circuit
* ============================================================================
* fc = R/(2*pi*L) = 1000/(2*pi*0.1) ≈ 1591.5 Hz
*
* Tests inductor WDF element.
* ============================================================================

L1 v_in v_out 100m
R1 v_out 0 1k
