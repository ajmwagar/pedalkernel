* ============================================================================
* Phase All-Pass Stage - Single JFET + Op-Amp
* PedalKernel Validation Circuit
* ============================================================================
* First-order all-pass filter for phaser circuits.
* JFET (2N5952) acts as voltage-controlled resistor in triode region.
* Op-amp provides unity-gain buffering.
* ============================================================================

* Supply
VCC vcc 0 DC 9

* Virtual ground (Vref = Vcc/2 = 4.5V)
R_vref1 vcc vref 470k
R_vref2 vref 0 470k
C_vref vref 0 10u

* Input coupling (AC couples to Vref bias)
C_in v_in vin_ac 100n
R_in vin_ac vref 1MEG

* All-pass network
* Standard first-order all-pass: R in series, RC to virtual ground via JFET
R_ap vin_ac vap 24k

* JFET as variable resistor (source follower config for Rds)
* Drain to ground, source is the resistive element
J1 0 vgate vap JMOD
C_ap vap vneg 47n

* JFET gate bias - divider from Vref
R_jb1 vref vgate 150k
R_jb2 vgate 0 150k

* Op-amp unity buffer (TL072)
* Uses simple VCVS model - we just need unity gain behavior
E_opamp vopout vref vneg vref 100k
R_opfb vneg vopout 100

* Output coupling
C_out vopout vout_ac 100n
R_load vout_ac 0 10k

* Output measurement
Eout v_out 0 vout_ac 0 1

* 2N5952 JFET model
.MODEL JMOD NJF(VTO=-4.0 BETA=0.5m LAMBDA=0.02 IS=1e-14 CGS=4p CGD=1.5p)
